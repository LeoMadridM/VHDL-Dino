--Melisa Saucedo Sánchez A01748077
--CONTADOR DE 10 BITS PARA CONTAR HASTA 525 DE LA VERTICAL DEL VGA 

----	CONTADOR A 524

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONT_V525 IS
	PORT(CLK, RESET : IN STD_LOGIC;
			ENA        : IN STD_LOGIC; 
			VSYNC      : OUT STD_LOGIC;
			COUNT      : OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END ENTITY;

ARCHITECTURE ARC OF CONT_V525 IS

	SIGNAL C1    : STD_LOGIC_VECTOR(9 DOWNTO 0);
	SIGNAL E, VS : STD_LOGIC;

 BEGIN	
	
	PR1 : PROCESS(CLK,RESET)
	
	BEGIN
		
		IF(RESET = '0') THEN
			C1 <= (OTHERS => '0');
		ELSIF (CLK'EVENT and CLK = '1' and ENA = '1') THEN
			IF C1 = "1000001100" THEN
				C1 <= (OTHERS => '0');
				
			ELSE
				C1 <= C1 + 1;
				
		   END IF;
		END IF;
	END PROCESS;
	
	COUNT <= C1;	
	
	PR2: PROCESS (C1)
	BEGIN
		IF (C1 > "0000000001") THEN
			VS <= '1';
		ELSE 
			VS <= '0';
		END IF;
	END PROCESS;
	
	VSYNC <= VS;	
		
END ARCHITECTURE;